----------------------------------------------------------------------------------
-- Company: UnB
-- Engineer: Rodrigo
-- 
-- Create Date: 17:12:09 05/31/2015 
-- Design Name: Rodrigo
-- Module Name: equ - Behavioral 
-- Project Name: Matrix Equation
----------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE work.dataTypes.ALL;

ENTITY equ IS
--	PORT (inputOne : IN STD_LOGIC_VECTOR (143 DOWNTO 0); -- 144 bits
--			inputTwo : IN STD_LOGIC_VECTOR (95 DOWNTO 0); -- 96 bits
--			operation : IN STD_LOGIC_VECTOR (2 DOWNTO 0); -- 3 bits
--			outputEQU : OUT STD_LOGIC_VECTOR (95 DOWNTO 0);
--			clkEQU : IN STD_LOGIC;
--			resetEQU : IN STD_LOGIC;
--			readyEQU : OUT STD_LOGIC
--			); -- 96 bits
END equ;

ARCHITECTURE Behavioral OF equ IS
BEGIN
END Behavioral;

